module MM(clk,i,j,reset,read,write,index,read_data,write_data,finish);

endmodule
